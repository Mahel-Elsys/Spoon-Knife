entity toto is (
  whatever : in std_logic;
  sig      : out std_logic );
end entity;
